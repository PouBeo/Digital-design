// File: FirPkg.sv
package FirPkg;
  parameter int WD_IN  = 24;
  parameter int WD_OUT = 24;
  parameter int DATA_WIDTH = 24;
  parameter int N_TAP = 32;

endpackage
